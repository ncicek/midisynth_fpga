`timescale 10ns / 10ns
module tuning_code_lookup(
	input wire [6:0] midi_byte,
	output reg [31:0] tuning_code
);

	always @* begin
		case(midi_byte)
			7'd0:	tuning_code = 32'd732;
			7'd1:	tuning_code = 32'd775;
			7'd2:	tuning_code = 32'd821;
			7'd3:	tuning_code = 32'd870;
			7'd4:	tuning_code = 32'd922;
			7'd5:	tuning_code = 32'd977;
			7'd6:	tuning_code = 32'd1035;
			7'd7:	tuning_code = 32'd1096;
			7'd8:	tuning_code = 32'd1161;
			7'd9:	tuning_code = 32'd1230;
			7'd10:	tuning_code = 32'd1303;
			7'd11:	tuning_code = 32'd1381;
			7'd12:	tuning_code = 32'd1463;
			7'd13:	tuning_code = 32'd1550;
			7'd14:	tuning_code = 32'd1642;
			7'd15:	tuning_code = 32'd1740;
			7'd16:	tuning_code = 32'd1843;
			7'd17:	tuning_code = 32'd1953;
			7'd18:	tuning_code = 32'd2069;
			7'd19:	tuning_code = 32'd2192;
			7'd20:	tuning_code = 32'd2323;
			7'd21:	tuning_code = 32'd2461;
			7'd22:	tuning_code = 32'd2607;
			7'd23:	tuning_code = 32'd2762;
			7'd24:	tuning_code = 32'd2926;
			7'd25:	tuning_code = 32'd3100;
			7'd26:	tuning_code = 32'd3285;
			7'd27:	tuning_code = 32'd3480;
			7'd28:	tuning_code = 32'd3687;
			7'd29:	tuning_code = 32'd3906;
			7'd30:	tuning_code = 32'd4138;
			7'd31:	tuning_code = 32'd4384;
			7'd32:	tuning_code = 32'd4645;
			7'd33:	tuning_code = 32'd4921;
			7'd34:	tuning_code = 32'd5214;
			7'd35:	tuning_code = 32'd5524;
			7'd36:	tuning_code = 32'd5852;
			7'd37:	tuning_code = 32'd6200;
			7'd38:	tuning_code = 32'd6569;
			7'd39:	tuning_code = 32'd6960;
			7'd40:	tuning_code = 32'd7374;
			7'd41:	tuning_code = 32'd7812;
			7'd42:	tuning_code = 32'd8277;
			7'd43:	tuning_code = 32'd8769;
			7'd44:	tuning_code = 32'd9290;
			7'd45:	tuning_code = 32'd9843;
			7'd46:	tuning_code = 32'd10428;
			7'd47:	tuning_code = 32'd11048;
			7'd48:	tuning_code = 32'd11705;
			7'd49:	tuning_code = 32'd12401;
			7'd50:	tuning_code = 32'd13138;
			7'd51:	tuning_code = 32'd13920;
			7'd52:	tuning_code = 32'd14747;
			7'd53:	tuning_code = 32'd15624;
			7'd54:	tuning_code = 32'd16553;
			7'd55:	tuning_code = 32'd17538;
			7'd56:	tuning_code = 32'd18580;
			7'd57:	tuning_code = 32'd19685;
			7'd58:	tuning_code = 32'd20856;
			7'd59:	tuning_code = 32'd22096;
			7'd60:	tuning_code = 32'd23410;
			7'd61:	tuning_code = 32'd24802;
			7'd62:	tuning_code = 32'd26277;
			7'd63:	tuning_code = 32'd27839;
			7'd64:	tuning_code = 32'd29495;
			7'd65:	tuning_code = 32'd31248;
			7'd66:	tuning_code = 32'd33107;
			7'd67:	tuning_code = 32'd35075;
			7'd68:	tuning_code = 32'd37161;
			7'd69:	tuning_code = 32'd39371;
			7'd70:	tuning_code = 32'd41712;
			7'd71:	tuning_code = 32'd44192;
			7'd72:	tuning_code = 32'd46820;
			7'd73:	tuning_code = 32'd49604;
			7'd74:	tuning_code = 32'd52553;
			7'd75:	tuning_code = 32'd55678;
			7'd76:	tuning_code = 32'd58989;
			7'd77:	tuning_code = 32'd62497;
			7'd78:	tuning_code = 32'd66213;
			7'd79:	tuning_code = 32'd70150;
			7'd80:	tuning_code = 32'd74322;
			7'd81:	tuning_code = 32'd78741;
			7'd82:	tuning_code = 32'd83423;
			7'd83:	tuning_code = 32'd88384;
			7'd84:	tuning_code = 32'd93639;
			7'd85:	tuning_code = 32'd99208;
			7'd86:	tuning_code = 32'd105107;
			7'd87:	tuning_code = 32'd111357;
			7'd88:	tuning_code = 32'd117978;
			7'd89:	tuning_code = 32'd124994;
			7'd90:	tuning_code = 32'd132426;
			7'd91:	tuning_code = 32'd140301;
			7'd92:	tuning_code = 32'd148643;
			7'd93:	tuning_code = 32'd157482;
			7'd94:	tuning_code = 32'd166847;
			7'd95:	tuning_code = 32'd176768;
			7'd96:	tuning_code = 32'd187279;
			7'd97:	tuning_code = 32'd198415;
			7'd98:	tuning_code = 32'd210213;
			7'd99:	tuning_code = 32'd222713;
			7'd100:	tuning_code = 32'd235957;
			7'd101:	tuning_code = 32'd249987;
			7'd102:	tuning_code = 32'd264852;
			7'd103:	tuning_code = 32'd280601;
			7'd104:	tuning_code = 32'd297287;
			7'd105:	tuning_code = 32'd314964;
			7'd106:	tuning_code = 32'd333693;
			7'd107:	tuning_code = 32'd353535;
			7'd108:	tuning_code = 32'd374558;
			7'd109:	tuning_code = 32'd396830;
			7'd110:	tuning_code = 32'd420427;
			7'd111:	tuning_code = 32'd445427;
			7'd112:	tuning_code = 32'd471913;
			7'd113:	tuning_code = 32'd499975;
			7'd114:	tuning_code = 32'd529705;
			7'd115:	tuning_code = 32'd561203;
			7'd116:	tuning_code = 32'd594573;
			7'd117:	tuning_code = 32'd629929;
			7'd118:	tuning_code = 32'd667386;
			7'd119:	tuning_code = 32'd707071;
			7'd120:	tuning_code = 32'd749115;
			7'd121:	tuning_code = 32'd793660;
			7'd122:	tuning_code = 32'd840854;
			7'd123:	tuning_code = 32'd890853;
			7'd124:	tuning_code = 32'd943826;
			7'd125:	tuning_code = 32'd999949;
			7'd126:	tuning_code = 32'd1059409;
			default: tuning_code = 32'd66213;
		endcase
	end
endmodule