module ram (din, addr, write_en, clk, dout);
  parameter addr_width = 8;
  parameter data_width = 8;
  input [addr_width-1:0] addr;
  input [data_width-1:0] din;
  input wire write_en;
  input wire clk;	  
  output wire [data_width-1:0] dout;
  reg [data_width-1:0] mem [(1<<addr_width)-1:0];
    // Define RAM as an indexed memory array.

  always @(posedge clk) // Control with a clock edge.
  begin
    if (write_en) // And control with a write enable.
      mem[(addr)] <= din;
  end
  assign dout = mem[addr];	  
  
  //initial 
//	  
//	begin
//		integer i;
//		for (i=0; i<100000; i=i+1) mem[i] <= 128'b0;
//	end
endmodule
