module sine_table(
	//input wire i_clk,
	input wire [9:0] theta,
	output reg signed [15:0] sine_sample
);

	always @(theta) begin
		case(theta)
			10'd0:	sine_sample = -16'sd0;
			10'd1:	sine_sample = -16'sd201;
			10'd2:	sine_sample = -16'sd402;
			10'd3:	sine_sample = -16'sd603;
			10'd4:	sine_sample = -16'sd804;
			10'd5:	sine_sample = -16'sd1005;
			10'd6:	sine_sample = -16'sd1206;
			10'd7:	sine_sample = -16'sd1407;
			10'd8:	sine_sample = -16'sd1608;
			10'd9:	sine_sample = -16'sd1809;
			10'd10:	sine_sample = -16'sd2009;
			10'd11:	sine_sample = -16'sd2210;
			10'd12:	sine_sample = -16'sd2411;
			10'd13:	sine_sample = -16'sd2611;
			10'd14:	sine_sample = -16'sd2811;
			10'd15:	sine_sample = -16'sd3012;
			10'd16:	sine_sample = -16'sd3212;
			10'd17:	sine_sample = -16'sd3412;
			10'd18:	sine_sample = -16'sd3612;
			10'd19:	sine_sample = -16'sd3812;
			10'd20:	sine_sample = -16'sd4011;
			10'd21:	sine_sample = -16'sd4211;
			10'd22:	sine_sample = -16'sd4410;
			10'd23:	sine_sample = -16'sd4609;
			10'd24:	sine_sample = -16'sd4808;
			10'd25:	sine_sample = -16'sd5007;
			10'd26:	sine_sample = -16'sd5205;
			10'd27:	sine_sample = -16'sd5404;
			10'd28:	sine_sample = -16'sd5602;
			10'd29:	sine_sample = -16'sd5800;
			10'd30:	sine_sample = -16'sd5998;
			10'd31:	sine_sample = -16'sd6195;
			10'd32:	sine_sample = -16'sd6393;
			10'd33:	sine_sample = -16'sd6590;
			10'd34:	sine_sample = -16'sd6787;
			10'd35:	sine_sample = -16'sd6983;
			10'd36:	sine_sample = -16'sd7180;
			10'd37:	sine_sample = -16'sd7376;
			10'd38:	sine_sample = -16'sd7571;
			10'd39:	sine_sample = -16'sd7767;
			10'd40:	sine_sample = -16'sd7962;
			10'd41:	sine_sample = -16'sd8157;
			10'd42:	sine_sample = -16'sd8351;
			10'd43:	sine_sample = -16'sd8546;
			10'd44:	sine_sample = -16'sd8740;
			10'd45:	sine_sample = -16'sd8933;
			10'd46:	sine_sample = -16'sd9127;
			10'd47:	sine_sample = -16'sd9319;
			10'd48:	sine_sample = -16'sd9512;
			10'd49:	sine_sample = -16'sd9704;
			10'd50:	sine_sample = -16'sd9896;
			10'd51:	sine_sample = -16'sd10088;
			10'd52:	sine_sample = -16'sd10279;
			10'd53:	sine_sample = -16'sd10469;
			10'd54:	sine_sample = -16'sd10660;
			10'd55:	sine_sample = -16'sd10850;
			10'd56:	sine_sample = -16'sd11039;
			10'd57:	sine_sample = -16'sd11228;
			10'd58:	sine_sample = -16'sd11417;
			10'd59:	sine_sample = -16'sd11605;
			10'd60:	sine_sample = -16'sd11793;
			10'd61:	sine_sample = -16'sd11980;
			10'd62:	sine_sample = -16'sd12167;
			10'd63:	sine_sample = -16'sd12354;
			10'd64:	sine_sample = -16'sd12540;
			10'd65:	sine_sample = -16'sd12725;
			10'd66:	sine_sample = -16'sd12910;
			10'd67:	sine_sample = -16'sd13095;
			10'd68:	sine_sample = -16'sd13279;
			10'd69:	sine_sample = -16'sd13463;
			10'd70:	sine_sample = -16'sd13646;
			10'd71:	sine_sample = -16'sd13828;
			10'd72:	sine_sample = -16'sd14010;
			10'd73:	sine_sample = -16'sd14192;
			10'd74:	sine_sample = -16'sd14373;
			10'd75:	sine_sample = -16'sd14553;
			10'd76:	sine_sample = -16'sd14733;
			10'd77:	sine_sample = -16'sd14912;
			10'd78:	sine_sample = -16'sd15091;
			10'd79:	sine_sample = -16'sd15269;
			10'd80:	sine_sample = -16'sd15447;
			10'd81:	sine_sample = -16'sd15624;
			10'd82:	sine_sample = -16'sd15800;
			10'd83:	sine_sample = -16'sd15976;
			10'd84:	sine_sample = -16'sd16151;
			10'd85:	sine_sample = -16'sd16326;
			10'd86:	sine_sample = -16'sd16500;
			10'd87:	sine_sample = -16'sd16673;
			10'd88:	sine_sample = -16'sd16846;
			10'd89:	sine_sample = -16'sd17018;
			10'd90:	sine_sample = -16'sd17190;
			10'd91:	sine_sample = -16'sd17361;
			10'd92:	sine_sample = -16'sd17531;
			10'd93:	sine_sample = -16'sd17700;
			10'd94:	sine_sample = -16'sd17869;
			10'd95:	sine_sample = -16'sd18037;
			10'd96:	sine_sample = -16'sd18205;
			10'd97:	sine_sample = -16'sd18372;
			10'd98:	sine_sample = -16'sd18538;
			10'd99:	sine_sample = -16'sd18703;
			10'd100:	sine_sample = -16'sd18868;
			10'd101:	sine_sample = -16'sd19032;
			10'd102:	sine_sample = -16'sd19195;
			10'd103:	sine_sample = -16'sd19358;
			10'd104:	sine_sample = -16'sd19520;
			10'd105:	sine_sample = -16'sd19681;
			10'd106:	sine_sample = -16'sd19841;
			10'd107:	sine_sample = -16'sd20001;
			10'd108:	sine_sample = -16'sd20160;
			10'd109:	sine_sample = -16'sd20318;
			10'd110:	sine_sample = -16'sd20475;
			10'd111:	sine_sample = -16'sd20632;
			10'd112:	sine_sample = -16'sd20788;
			10'd113:	sine_sample = -16'sd20943;
			10'd114:	sine_sample = -16'sd21097;
			10'd115:	sine_sample = -16'sd21251;
			10'd116:	sine_sample = -16'sd21403;
			10'd117:	sine_sample = -16'sd21555;
			10'd118:	sine_sample = -16'sd21706;
			10'd119:	sine_sample = -16'sd21856;
			10'd120:	sine_sample = -16'sd22006;
			10'd121:	sine_sample = -16'sd22154;
			10'd122:	sine_sample = -16'sd22302;
			10'd123:	sine_sample = -16'sd22449;
			10'd124:	sine_sample = -16'sd22595;
			10'd125:	sine_sample = -16'sd22740;
			10'd126:	sine_sample = -16'sd22884;
			10'd127:	sine_sample = -16'sd23028;
			10'd128:	sine_sample = -16'sd23170;
			10'd129:	sine_sample = -16'sd23312;
			10'd130:	sine_sample = -16'sd23453;
			10'd131:	sine_sample = -16'sd23593;
			10'd132:	sine_sample = -16'sd23732;
			10'd133:	sine_sample = -16'sd23870;
			10'd134:	sine_sample = -16'sd24008;
			10'd135:	sine_sample = -16'sd24144;
			10'd136:	sine_sample = -16'sd24279;
			10'd137:	sine_sample = -16'sd24414;
			10'd138:	sine_sample = -16'sd24548;
			10'd139:	sine_sample = -16'sd24680;
			10'd140:	sine_sample = -16'sd24812;
			10'd141:	sine_sample = -16'sd24943;
			10'd142:	sine_sample = -16'sd25073;
			10'd143:	sine_sample = -16'sd25202;
			10'd144:	sine_sample = -16'sd25330;
			10'd145:	sine_sample = -16'sd25457;
			10'd146:	sine_sample = -16'sd25583;
			10'd147:	sine_sample = -16'sd25708;
			10'd148:	sine_sample = -16'sd25833;
			10'd149:	sine_sample = -16'sd25956;
			10'd150:	sine_sample = -16'sd26078;
			10'd151:	sine_sample = -16'sd26199;
			10'd152:	sine_sample = -16'sd26320;
			10'd153:	sine_sample = -16'sd26439;
			10'd154:	sine_sample = -16'sd26557;
			10'd155:	sine_sample = -16'sd26674;
			10'd156:	sine_sample = -16'sd26791;
			10'd157:	sine_sample = -16'sd26906;
			10'd158:	sine_sample = -16'sd27020;
			10'd159:	sine_sample = -16'sd27133;
			10'd160:	sine_sample = -16'sd27246;
			10'd161:	sine_sample = -16'sd27357;
			10'd162:	sine_sample = -16'sd27467;
			10'd163:	sine_sample = -16'sd27576;
			10'd164:	sine_sample = -16'sd27684;
			10'd165:	sine_sample = -16'sd27791;
			10'd166:	sine_sample = -16'sd27897;
			10'd167:	sine_sample = -16'sd28002;
			10'd168:	sine_sample = -16'sd28106;
			10'd169:	sine_sample = -16'sd28209;
			10'd170:	sine_sample = -16'sd28311;
			10'd171:	sine_sample = -16'sd28411;
			10'd172:	sine_sample = -16'sd28511;
			10'd173:	sine_sample = -16'sd28610;
			10'd174:	sine_sample = -16'sd28707;
			10'd175:	sine_sample = -16'sd28803;
			10'd176:	sine_sample = -16'sd28899;
			10'd177:	sine_sample = -16'sd28993;
			10'd178:	sine_sample = -16'sd29086;
			10'd179:	sine_sample = -16'sd29178;
			10'd180:	sine_sample = -16'sd29269;
			10'd181:	sine_sample = -16'sd29359;
			10'd182:	sine_sample = -16'sd29448;
			10'd183:	sine_sample = -16'sd29535;
			10'd184:	sine_sample = -16'sd29622;
			10'd185:	sine_sample = -16'sd29707;
			10'd186:	sine_sample = -16'sd29792;
			10'd187:	sine_sample = -16'sd29875;
			10'd188:	sine_sample = -16'sd29957;
			10'd189:	sine_sample = -16'sd30038;
			10'd190:	sine_sample = -16'sd30118;
			10'd191:	sine_sample = -16'sd30196;
			10'd192:	sine_sample = -16'sd30274;
			10'd193:	sine_sample = -16'sd30350;
			10'd194:	sine_sample = -16'sd30425;
			10'd195:	sine_sample = -16'sd30499;
			10'd196:	sine_sample = -16'sd30572;
			10'd197:	sine_sample = -16'sd30644;
			10'd198:	sine_sample = -16'sd30715;
			10'd199:	sine_sample = -16'sd30784;
			10'd200:	sine_sample = -16'sd30853;
			10'd201:	sine_sample = -16'sd30920;
			10'd202:	sine_sample = -16'sd30986;
			10'd203:	sine_sample = -16'sd31050;
			10'd204:	sine_sample = -16'sd31114;
			10'd205:	sine_sample = -16'sd31177;
			10'd206:	sine_sample = -16'sd31238;
			10'd207:	sine_sample = -16'sd31298;
			10'd208:	sine_sample = -16'sd31357;
			10'd209:	sine_sample = -16'sd31415;
			10'd210:	sine_sample = -16'sd31471;
			10'd211:	sine_sample = -16'sd31527;
			10'd212:	sine_sample = -16'sd31581;
			10'd213:	sine_sample = -16'sd31634;
			10'd214:	sine_sample = -16'sd31686;
			10'd215:	sine_sample = -16'sd31737;
			10'd216:	sine_sample = -16'sd31786;
			10'd217:	sine_sample = -16'sd31834;
			10'd218:	sine_sample = -16'sd31881;
			10'd219:	sine_sample = -16'sd31927;
			10'd220:	sine_sample = -16'sd31972;
			10'd221:	sine_sample = -16'sd32015;
			10'd222:	sine_sample = -16'sd32058;
			10'd223:	sine_sample = -16'sd32099;
			10'd224:	sine_sample = -16'sd32138;
			10'd225:	sine_sample = -16'sd32177;
			10'd226:	sine_sample = -16'sd32214;
			10'd227:	sine_sample = -16'sd32251;
			10'd228:	sine_sample = -16'sd32286;
			10'd229:	sine_sample = -16'sd32319;
			10'd230:	sine_sample = -16'sd32352;
			10'd231:	sine_sample = -16'sd32383;
			10'd232:	sine_sample = -16'sd32413;
			10'd233:	sine_sample = -16'sd32442;
			10'd234:	sine_sample = -16'sd32470;
			10'd235:	sine_sample = -16'sd32496;
			10'd236:	sine_sample = -16'sd32522;
			10'd237:	sine_sample = -16'sd32546;
			10'd238:	sine_sample = -16'sd32568;
			10'd239:	sine_sample = -16'sd32590;
			10'd240:	sine_sample = -16'sd32610;
			10'd241:	sine_sample = -16'sd32629;
			10'd242:	sine_sample = -16'sd32647;
			10'd243:	sine_sample = -16'sd32664;
			10'd244:	sine_sample = -16'sd32679;
			10'd245:	sine_sample = -16'sd32693;
			10'd246:	sine_sample = -16'sd32706;
			10'd247:	sine_sample = -16'sd32718;
			10'd248:	sine_sample = -16'sd32729;
			10'd249:	sine_sample = -16'sd32738;
			10'd250:	sine_sample = -16'sd32746;
			10'd251:	sine_sample = -16'sd32753;
			10'd252:	sine_sample = -16'sd32758;
			10'd253:	sine_sample = -16'sd32762;
			10'd254:	sine_sample = -16'sd32766;
			10'd255:	sine_sample = -16'sd32767;
			10'd256:	sine_sample = -16'sd32768;
			10'd257:	sine_sample = -16'sd32767;
			10'd258:	sine_sample = -16'sd32766;
			10'd259:	sine_sample = -16'sd32762;
			10'd260:	sine_sample = -16'sd32758;
			10'd261:	sine_sample = -16'sd32753;
			10'd262:	sine_sample = -16'sd32746;
			10'd263:	sine_sample = -16'sd32738;
			10'd264:	sine_sample = -16'sd32729;
			10'd265:	sine_sample = -16'sd32718;
			10'd266:	sine_sample = -16'sd32706;
			10'd267:	sine_sample = -16'sd32693;
			10'd268:	sine_sample = -16'sd32679;
			10'd269:	sine_sample = -16'sd32664;
			10'd270:	sine_sample = -16'sd32647;
			10'd271:	sine_sample = -16'sd32629;
			10'd272:	sine_sample = -16'sd32610;
			10'd273:	sine_sample = -16'sd32590;
			10'd274:	sine_sample = -16'sd32568;
			10'd275:	sine_sample = -16'sd32546;
			10'd276:	sine_sample = -16'sd32522;
			10'd277:	sine_sample = -16'sd32496;
			10'd278:	sine_sample = -16'sd32470;
			10'd279:	sine_sample = -16'sd32442;
			10'd280:	sine_sample = -16'sd32413;
			10'd281:	sine_sample = -16'sd32383;
			10'd282:	sine_sample = -16'sd32352;
			10'd283:	sine_sample = -16'sd32319;
			10'd284:	sine_sample = -16'sd32286;
			10'd285:	sine_sample = -16'sd32251;
			10'd286:	sine_sample = -16'sd32214;
			10'd287:	sine_sample = -16'sd32177;
			10'd288:	sine_sample = -16'sd32138;
			10'd289:	sine_sample = -16'sd32099;
			10'd290:	sine_sample = -16'sd32058;
			10'd291:	sine_sample = -16'sd32015;
			10'd292:	sine_sample = -16'sd31972;
			10'd293:	sine_sample = -16'sd31927;
			10'd294:	sine_sample = -16'sd31881;
			10'd295:	sine_sample = -16'sd31834;
			10'd296:	sine_sample = -16'sd31786;
			10'd297:	sine_sample = -16'sd31737;
			10'd298:	sine_sample = -16'sd31686;
			10'd299:	sine_sample = -16'sd31634;
			10'd300:	sine_sample = -16'sd31581;
			10'd301:	sine_sample = -16'sd31527;
			10'd302:	sine_sample = -16'sd31471;
			10'd303:	sine_sample = -16'sd31415;
			10'd304:	sine_sample = -16'sd31357;
			10'd305:	sine_sample = -16'sd31298;
			10'd306:	sine_sample = -16'sd31238;
			10'd307:	sine_sample = -16'sd31177;
			10'd308:	sine_sample = -16'sd31114;
			10'd309:	sine_sample = -16'sd31050;
			10'd310:	sine_sample = -16'sd30986;
			10'd311:	sine_sample = -16'sd30920;
			10'd312:	sine_sample = -16'sd30853;
			10'd313:	sine_sample = -16'sd30784;
			10'd314:	sine_sample = -16'sd30715;
			10'd315:	sine_sample = -16'sd30644;
			10'd316:	sine_sample = -16'sd30572;
			10'd317:	sine_sample = -16'sd30499;
			10'd318:	sine_sample = -16'sd30425;
			10'd319:	sine_sample = -16'sd30350;
			10'd320:	sine_sample = -16'sd30274;
			10'd321:	sine_sample = -16'sd30196;
			10'd322:	sine_sample = -16'sd30118;
			10'd323:	sine_sample = -16'sd30038;
			10'd324:	sine_sample = -16'sd29957;
			10'd325:	sine_sample = -16'sd29875;
			10'd326:	sine_sample = -16'sd29792;
			10'd327:	sine_sample = -16'sd29707;
			10'd328:	sine_sample = -16'sd29622;
			10'd329:	sine_sample = -16'sd29535;
			10'd330:	sine_sample = -16'sd29448;
			10'd331:	sine_sample = -16'sd29359;
			10'd332:	sine_sample = -16'sd29269;
			10'd333:	sine_sample = -16'sd29178;
			10'd334:	sine_sample = -16'sd29086;
			10'd335:	sine_sample = -16'sd28993;
			10'd336:	sine_sample = -16'sd28899;
			10'd337:	sine_sample = -16'sd28803;
			10'd338:	sine_sample = -16'sd28707;
			10'd339:	sine_sample = -16'sd28610;
			10'd340:	sine_sample = -16'sd28511;
			10'd341:	sine_sample = -16'sd28411;
			10'd342:	sine_sample = -16'sd28311;
			10'd343:	sine_sample = -16'sd28209;
			10'd344:	sine_sample = -16'sd28106;
			10'd345:	sine_sample = -16'sd28002;
			10'd346:	sine_sample = -16'sd27897;
			10'd347:	sine_sample = -16'sd27791;
			10'd348:	sine_sample = -16'sd27684;
			10'd349:	sine_sample = -16'sd27576;
			10'd350:	sine_sample = -16'sd27467;
			10'd351:	sine_sample = -16'sd27357;
			10'd352:	sine_sample = -16'sd27246;
			10'd353:	sine_sample = -16'sd27133;
			10'd354:	sine_sample = -16'sd27020;
			10'd355:	sine_sample = -16'sd26906;
			10'd356:	sine_sample = -16'sd26791;
			10'd357:	sine_sample = -16'sd26674;
			10'd358:	sine_sample = -16'sd26557;
			10'd359:	sine_sample = -16'sd26439;
			10'd360:	sine_sample = -16'sd26320;
			10'd361:	sine_sample = -16'sd26199;
			10'd362:	sine_sample = -16'sd26078;
			10'd363:	sine_sample = -16'sd25956;
			10'd364:	sine_sample = -16'sd25833;
			10'd365:	sine_sample = -16'sd25708;
			10'd366:	sine_sample = -16'sd25583;
			10'd367:	sine_sample = -16'sd25457;
			10'd368:	sine_sample = -16'sd25330;
			10'd369:	sine_sample = -16'sd25202;
			10'd370:	sine_sample = -16'sd25073;
			10'd371:	sine_sample = -16'sd24943;
			10'd372:	sine_sample = -16'sd24812;
			10'd373:	sine_sample = -16'sd24680;
			10'd374:	sine_sample = -16'sd24548;
			10'd375:	sine_sample = -16'sd24414;
			10'd376:	sine_sample = -16'sd24279;
			10'd377:	sine_sample = -16'sd24144;
			10'd378:	sine_sample = -16'sd24008;
			10'd379:	sine_sample = -16'sd23870;
			10'd380:	sine_sample = -16'sd23732;
			10'd381:	sine_sample = -16'sd23593;
			10'd382:	sine_sample = -16'sd23453;
			10'd383:	sine_sample = -16'sd23312;
			10'd384:	sine_sample = -16'sd23170;
			10'd385:	sine_sample = -16'sd23028;
			10'd386:	sine_sample = -16'sd22884;
			10'd387:	sine_sample = -16'sd22740;
			10'd388:	sine_sample = -16'sd22595;
			10'd389:	sine_sample = -16'sd22449;
			10'd390:	sine_sample = -16'sd22302;
			10'd391:	sine_sample = -16'sd22154;
			10'd392:	sine_sample = -16'sd22006;
			10'd393:	sine_sample = -16'sd21856;
			10'd394:	sine_sample = -16'sd21706;
			10'd395:	sine_sample = -16'sd21555;
			10'd396:	sine_sample = -16'sd21403;
			10'd397:	sine_sample = -16'sd21251;
			10'd398:	sine_sample = -16'sd21097;
			10'd399:	sine_sample = -16'sd20943;
			10'd400:	sine_sample = -16'sd20788;
			10'd401:	sine_sample = -16'sd20632;
			10'd402:	sine_sample = -16'sd20475;
			10'd403:	sine_sample = -16'sd20318;
			10'd404:	sine_sample = -16'sd20160;
			10'd405:	sine_sample = -16'sd20001;
			10'd406:	sine_sample = -16'sd19841;
			10'd407:	sine_sample = -16'sd19681;
			10'd408:	sine_sample = -16'sd19520;
			10'd409:	sine_sample = -16'sd19358;
			10'd410:	sine_sample = -16'sd19195;
			10'd411:	sine_sample = -16'sd19032;
			10'd412:	sine_sample = -16'sd18868;
			10'd413:	sine_sample = -16'sd18703;
			10'd414:	sine_sample = -16'sd18538;
			10'd415:	sine_sample = -16'sd18372;
			10'd416:	sine_sample = -16'sd18205;
			10'd417:	sine_sample = -16'sd18037;
			10'd418:	sine_sample = -16'sd17869;
			10'd419:	sine_sample = -16'sd17700;
			10'd420:	sine_sample = -16'sd17531;
			10'd421:	sine_sample = -16'sd17361;
			10'd422:	sine_sample = -16'sd17190;
			10'd423:	sine_sample = -16'sd17018;
			10'd424:	sine_sample = -16'sd16846;
			10'd425:	sine_sample = -16'sd16673;
			10'd426:	sine_sample = -16'sd16500;
			10'd427:	sine_sample = -16'sd16326;
			10'd428:	sine_sample = -16'sd16151;
			10'd429:	sine_sample = -16'sd15976;
			10'd430:	sine_sample = -16'sd15800;
			10'd431:	sine_sample = -16'sd15624;
			10'd432:	sine_sample = -16'sd15447;
			10'd433:	sine_sample = -16'sd15269;
			10'd434:	sine_sample = -16'sd15091;
			10'd435:	sine_sample = -16'sd14912;
			10'd436:	sine_sample = -16'sd14733;
			10'd437:	sine_sample = -16'sd14553;
			10'd438:	sine_sample = -16'sd14373;
			10'd439:	sine_sample = -16'sd14192;
			10'd440:	sine_sample = -16'sd14010;
			10'd441:	sine_sample = -16'sd13828;
			10'd442:	sine_sample = -16'sd13646;
			10'd443:	sine_sample = -16'sd13463;
			10'd444:	sine_sample = -16'sd13279;
			10'd445:	sine_sample = -16'sd13095;
			10'd446:	sine_sample = -16'sd12910;
			10'd447:	sine_sample = -16'sd12725;
			10'd448:	sine_sample = -16'sd12540;
			10'd449:	sine_sample = -16'sd12354;
			10'd450:	sine_sample = -16'sd12167;
			10'd451:	sine_sample = -16'sd11980;
			10'd452:	sine_sample = -16'sd11793;
			10'd453:	sine_sample = -16'sd11605;
			10'd454:	sine_sample = -16'sd11417;
			10'd455:	sine_sample = -16'sd11228;
			10'd456:	sine_sample = -16'sd11039;
			10'd457:	sine_sample = -16'sd10850;
			10'd458:	sine_sample = -16'sd10660;
			10'd459:	sine_sample = -16'sd10469;
			10'd460:	sine_sample = -16'sd10279;
			10'd461:	sine_sample = -16'sd10088;
			10'd462:	sine_sample = -16'sd9896;
			10'd463:	sine_sample = -16'sd9704;
			10'd464:	sine_sample = -16'sd9512;
			10'd465:	sine_sample = -16'sd9319;
			10'd466:	sine_sample = -16'sd9127;
			10'd467:	sine_sample = -16'sd8933;
			10'd468:	sine_sample = -16'sd8740;
			10'd469:	sine_sample = -16'sd8546;
			10'd470:	sine_sample = -16'sd8351;
			10'd471:	sine_sample = -16'sd8157;
			10'd472:	sine_sample = -16'sd7962;
			10'd473:	sine_sample = -16'sd7767;
			10'd474:	sine_sample = -16'sd7571;
			10'd475:	sine_sample = -16'sd7376;
			10'd476:	sine_sample = -16'sd7180;
			10'd477:	sine_sample = -16'sd6983;
			10'd478:	sine_sample = -16'sd6787;
			10'd479:	sine_sample = -16'sd6590;
			10'd480:	sine_sample = -16'sd6393;
			10'd481:	sine_sample = -16'sd6195;
			10'd482:	sine_sample = -16'sd5998;
			10'd483:	sine_sample = -16'sd5800;
			10'd484:	sine_sample = -16'sd5602;
			10'd485:	sine_sample = -16'sd5404;
			10'd486:	sine_sample = -16'sd5205;
			10'd487:	sine_sample = -16'sd5007;
			10'd488:	sine_sample = -16'sd4808;
			10'd489:	sine_sample = -16'sd4609;
			10'd490:	sine_sample = -16'sd4410;
			10'd491:	sine_sample = -16'sd4211;
			10'd492:	sine_sample = -16'sd4011;
			10'd493:	sine_sample = -16'sd3812;
			10'd494:	sine_sample = -16'sd3612;
			10'd495:	sine_sample = -16'sd3412;
			10'd496:	sine_sample = -16'sd3212;
			10'd497:	sine_sample = -16'sd3012;
			10'd498:	sine_sample = -16'sd2811;
			10'd499:	sine_sample = -16'sd2611;
			10'd500:	sine_sample = -16'sd2411;
			10'd501:	sine_sample = -16'sd2210;
			10'd502:	sine_sample = -16'sd2009;
			10'd503:	sine_sample = -16'sd1809;
			10'd504:	sine_sample = -16'sd1608;
			10'd505:	sine_sample = -16'sd1407;
			10'd506:	sine_sample = -16'sd1206;
			10'd507:	sine_sample = -16'sd1005;
			10'd508:	sine_sample = -16'sd804;
			10'd509:	sine_sample = -16'sd603;
			10'd510:	sine_sample = -16'sd402;
			10'd511:	sine_sample = -16'sd201;
			10'd512:	sine_sample = -16'sd0;
			10'd513:	sine_sample = 16'sd201;
			10'd514:	sine_sample = 16'sd402;
			10'd515:	sine_sample = 16'sd603;
			10'd516:	sine_sample = 16'sd804;
			10'd517:	sine_sample = 16'sd1005;
			10'd518:	sine_sample = 16'sd1206;
			10'd519:	sine_sample = 16'sd1407;
			10'd520:	sine_sample = 16'sd1608;
			10'd521:	sine_sample = 16'sd1809;
			10'd522:	sine_sample = 16'sd2009;
			10'd523:	sine_sample = 16'sd2210;
			10'd524:	sine_sample = 16'sd2411;
			10'd525:	sine_sample = 16'sd2611;
			10'd526:	sine_sample = 16'sd2811;
			10'd527:	sine_sample = 16'sd3012;
			10'd528:	sine_sample = 16'sd3212;
			10'd529:	sine_sample = 16'sd3412;
			10'd530:	sine_sample = 16'sd3612;
			10'd531:	sine_sample = 16'sd3812;
			10'd532:	sine_sample = 16'sd4011;
			10'd533:	sine_sample = 16'sd4211;
			10'd534:	sine_sample = 16'sd4410;
			10'd535:	sine_sample = 16'sd4609;
			10'd536:	sine_sample = 16'sd4808;
			10'd537:	sine_sample = 16'sd5007;
			10'd538:	sine_sample = 16'sd5205;
			10'd539:	sine_sample = 16'sd5404;
			10'd540:	sine_sample = 16'sd5602;
			10'd541:	sine_sample = 16'sd5800;
			10'd542:	sine_sample = 16'sd5998;
			10'd543:	sine_sample = 16'sd6195;
			10'd544:	sine_sample = 16'sd6393;
			10'd545:	sine_sample = 16'sd6590;
			10'd546:	sine_sample = 16'sd6787;
			10'd547:	sine_sample = 16'sd6983;
			10'd548:	sine_sample = 16'sd7180;
			10'd549:	sine_sample = 16'sd7376;
			10'd550:	sine_sample = 16'sd7571;
			10'd551:	sine_sample = 16'sd7767;
			10'd552:	sine_sample = 16'sd7962;
			10'd553:	sine_sample = 16'sd8157;
			10'd554:	sine_sample = 16'sd8351;
			10'd555:	sine_sample = 16'sd8546;
			10'd556:	sine_sample = 16'sd8740;
			10'd557:	sine_sample = 16'sd8933;
			10'd558:	sine_sample = 16'sd9127;
			10'd559:	sine_sample = 16'sd9319;
			10'd560:	sine_sample = 16'sd9512;
			10'd561:	sine_sample = 16'sd9704;
			10'd562:	sine_sample = 16'sd9896;
			10'd563:	sine_sample = 16'sd10088;
			10'd564:	sine_sample = 16'sd10279;
			10'd565:	sine_sample = 16'sd10469;
			10'd566:	sine_sample = 16'sd10660;
			10'd567:	sine_sample = 16'sd10850;
			10'd568:	sine_sample = 16'sd11039;
			10'd569:	sine_sample = 16'sd11228;
			10'd570:	sine_sample = 16'sd11417;
			10'd571:	sine_sample = 16'sd11605;
			10'd572:	sine_sample = 16'sd11793;
			10'd573:	sine_sample = 16'sd11980;
			10'd574:	sine_sample = 16'sd12167;
			10'd575:	sine_sample = 16'sd12354;
			10'd576:	sine_sample = 16'sd12540;
			10'd577:	sine_sample = 16'sd12725;
			10'd578:	sine_sample = 16'sd12910;
			10'd579:	sine_sample = 16'sd13095;
			10'd580:	sine_sample = 16'sd13279;
			10'd581:	sine_sample = 16'sd13463;
			10'd582:	sine_sample = 16'sd13646;
			10'd583:	sine_sample = 16'sd13828;
			10'd584:	sine_sample = 16'sd14010;
			10'd585:	sine_sample = 16'sd14192;
			10'd586:	sine_sample = 16'sd14373;
			10'd587:	sine_sample = 16'sd14553;
			10'd588:	sine_sample = 16'sd14733;
			10'd589:	sine_sample = 16'sd14912;
			10'd590:	sine_sample = 16'sd15091;
			10'd591:	sine_sample = 16'sd15269;
			10'd592:	sine_sample = 16'sd15447;
			10'd593:	sine_sample = 16'sd15624;
			10'd594:	sine_sample = 16'sd15800;
			10'd595:	sine_sample = 16'sd15976;
			10'd596:	sine_sample = 16'sd16151;
			10'd597:	sine_sample = 16'sd16326;
			10'd598:	sine_sample = 16'sd16500;
			10'd599:	sine_sample = 16'sd16673;
			10'd600:	sine_sample = 16'sd16846;
			10'd601:	sine_sample = 16'sd17018;
			10'd602:	sine_sample = 16'sd17190;
			10'd603:	sine_sample = 16'sd17361;
			10'd604:	sine_sample = 16'sd17531;
			10'd605:	sine_sample = 16'sd17700;
			10'd606:	sine_sample = 16'sd17869;
			10'd607:	sine_sample = 16'sd18037;
			10'd608:	sine_sample = 16'sd18205;
			10'd609:	sine_sample = 16'sd18372;
			10'd610:	sine_sample = 16'sd18538;
			10'd611:	sine_sample = 16'sd18703;
			10'd612:	sine_sample = 16'sd18868;
			10'd613:	sine_sample = 16'sd19032;
			10'd614:	sine_sample = 16'sd19195;
			10'd615:	sine_sample = 16'sd19358;
			10'd616:	sine_sample = 16'sd19520;
			10'd617:	sine_sample = 16'sd19681;
			10'd618:	sine_sample = 16'sd19841;
			10'd619:	sine_sample = 16'sd20001;
			10'd620:	sine_sample = 16'sd20160;
			10'd621:	sine_sample = 16'sd20318;
			10'd622:	sine_sample = 16'sd20475;
			10'd623:	sine_sample = 16'sd20632;
			10'd624:	sine_sample = 16'sd20788;
			10'd625:	sine_sample = 16'sd20943;
			10'd626:	sine_sample = 16'sd21097;
			10'd627:	sine_sample = 16'sd21251;
			10'd628:	sine_sample = 16'sd21403;
			10'd629:	sine_sample = 16'sd21555;
			10'd630:	sine_sample = 16'sd21706;
			10'd631:	sine_sample = 16'sd21856;
			10'd632:	sine_sample = 16'sd22006;
			10'd633:	sine_sample = 16'sd22154;
			10'd634:	sine_sample = 16'sd22302;
			10'd635:	sine_sample = 16'sd22449;
			10'd636:	sine_sample = 16'sd22595;
			10'd637:	sine_sample = 16'sd22740;
			10'd638:	sine_sample = 16'sd22884;
			10'd639:	sine_sample = 16'sd23028;
			10'd640:	sine_sample = 16'sd23170;
			10'd641:	sine_sample = 16'sd23312;
			10'd642:	sine_sample = 16'sd23453;
			10'd643:	sine_sample = 16'sd23593;
			10'd644:	sine_sample = 16'sd23732;
			10'd645:	sine_sample = 16'sd23870;
			10'd646:	sine_sample = 16'sd24008;
			10'd647:	sine_sample = 16'sd24144;
			10'd648:	sine_sample = 16'sd24279;
			10'd649:	sine_sample = 16'sd24414;
			10'd650:	sine_sample = 16'sd24548;
			10'd651:	sine_sample = 16'sd24680;
			10'd652:	sine_sample = 16'sd24812;
			10'd653:	sine_sample = 16'sd24943;
			10'd654:	sine_sample = 16'sd25073;
			10'd655:	sine_sample = 16'sd25202;
			10'd656:	sine_sample = 16'sd25330;
			10'd657:	sine_sample = 16'sd25457;
			10'd658:	sine_sample = 16'sd25583;
			10'd659:	sine_sample = 16'sd25708;
			10'd660:	sine_sample = 16'sd25833;
			10'd661:	sine_sample = 16'sd25956;
			10'd662:	sine_sample = 16'sd26078;
			10'd663:	sine_sample = 16'sd26199;
			10'd664:	sine_sample = 16'sd26320;
			10'd665:	sine_sample = 16'sd26439;
			10'd666:	sine_sample = 16'sd26557;
			10'd667:	sine_sample = 16'sd26674;
			10'd668:	sine_sample = 16'sd26791;
			10'd669:	sine_sample = 16'sd26906;
			10'd670:	sine_sample = 16'sd27020;
			10'd671:	sine_sample = 16'sd27133;
			10'd672:	sine_sample = 16'sd27246;
			10'd673:	sine_sample = 16'sd27357;
			10'd674:	sine_sample = 16'sd27467;
			10'd675:	sine_sample = 16'sd27576;
			10'd676:	sine_sample = 16'sd27684;
			10'd677:	sine_sample = 16'sd27791;
			10'd678:	sine_sample = 16'sd27897;
			10'd679:	sine_sample = 16'sd28002;
			10'd680:	sine_sample = 16'sd28106;
			10'd681:	sine_sample = 16'sd28209;
			10'd682:	sine_sample = 16'sd28311;
			10'd683:	sine_sample = 16'sd28411;
			10'd684:	sine_sample = 16'sd28511;
			10'd685:	sine_sample = 16'sd28610;
			10'd686:	sine_sample = 16'sd28707;
			10'd687:	sine_sample = 16'sd28803;
			10'd688:	sine_sample = 16'sd28899;
			10'd689:	sine_sample = 16'sd28993;
			10'd690:	sine_sample = 16'sd29086;
			10'd691:	sine_sample = 16'sd29178;
			10'd692:	sine_sample = 16'sd29269;
			10'd693:	sine_sample = 16'sd29359;
			10'd694:	sine_sample = 16'sd29448;
			10'd695:	sine_sample = 16'sd29535;
			10'd696:	sine_sample = 16'sd29622;
			10'd697:	sine_sample = 16'sd29707;
			10'd698:	sine_sample = 16'sd29792;
			10'd699:	sine_sample = 16'sd29875;
			10'd700:	sine_sample = 16'sd29957;
			10'd701:	sine_sample = 16'sd30038;
			10'd702:	sine_sample = 16'sd30118;
			10'd703:	sine_sample = 16'sd30196;
			10'd704:	sine_sample = 16'sd30274;
			10'd705:	sine_sample = 16'sd30350;
			10'd706:	sine_sample = 16'sd30425;
			10'd707:	sine_sample = 16'sd30499;
			10'd708:	sine_sample = 16'sd30572;
			10'd709:	sine_sample = 16'sd30644;
			10'd710:	sine_sample = 16'sd30715;
			10'd711:	sine_sample = 16'sd30784;
			10'd712:	sine_sample = 16'sd30853;
			10'd713:	sine_sample = 16'sd30920;
			10'd714:	sine_sample = 16'sd30986;
			10'd715:	sine_sample = 16'sd31050;
			10'd716:	sine_sample = 16'sd31114;
			10'd717:	sine_sample = 16'sd31177;
			10'd718:	sine_sample = 16'sd31238;
			10'd719:	sine_sample = 16'sd31298;
			10'd720:	sine_sample = 16'sd31357;
			10'd721:	sine_sample = 16'sd31415;
			10'd722:	sine_sample = 16'sd31471;
			10'd723:	sine_sample = 16'sd31527;
			10'd724:	sine_sample = 16'sd31581;
			10'd725:	sine_sample = 16'sd31634;
			10'd726:	sine_sample = 16'sd31686;
			10'd727:	sine_sample = 16'sd31737;
			10'd728:	sine_sample = 16'sd31786;
			10'd729:	sine_sample = 16'sd31834;
			10'd730:	sine_sample = 16'sd31881;
			10'd731:	sine_sample = 16'sd31927;
			10'd732:	sine_sample = 16'sd31972;
			10'd733:	sine_sample = 16'sd32015;
			10'd734:	sine_sample = 16'sd32058;
			10'd735:	sine_sample = 16'sd32099;
			10'd736:	sine_sample = 16'sd32138;
			10'd737:	sine_sample = 16'sd32177;
			10'd738:	sine_sample = 16'sd32214;
			10'd739:	sine_sample = 16'sd32251;
			10'd740:	sine_sample = 16'sd32286;
			10'd741:	sine_sample = 16'sd32319;
			10'd742:	sine_sample = 16'sd32352;
			10'd743:	sine_sample = 16'sd32383;
			10'd744:	sine_sample = 16'sd32413;
			10'd745:	sine_sample = 16'sd32442;
			10'd746:	sine_sample = 16'sd32470;
			10'd747:	sine_sample = 16'sd32496;
			10'd748:	sine_sample = 16'sd32522;
			10'd749:	sine_sample = 16'sd32546;
			10'd750:	sine_sample = 16'sd32568;
			10'd751:	sine_sample = 16'sd32590;
			10'd752:	sine_sample = 16'sd32610;
			10'd753:	sine_sample = 16'sd32629;
			10'd754:	sine_sample = 16'sd32647;
			10'd755:	sine_sample = 16'sd32664;
			10'd756:	sine_sample = 16'sd32679;
			10'd757:	sine_sample = 16'sd32693;
			10'd758:	sine_sample = 16'sd32706;
			10'd759:	sine_sample = 16'sd32718;
			10'd760:	sine_sample = 16'sd32729;
			10'd761:	sine_sample = 16'sd32738;
			10'd762:	sine_sample = 16'sd32746;
			10'd763:	sine_sample = 16'sd32753;
			10'd764:	sine_sample = 16'sd32758;
			10'd765:	sine_sample = 16'sd32762;
			10'd766:	sine_sample = 16'sd32766;
			10'd767:	sine_sample = 16'sd32767;
			10'd768:	sine_sample = 16'sd32768;
			10'd769:	sine_sample = 16'sd32767;
			10'd770:	sine_sample = 16'sd32766;
			10'd771:	sine_sample = 16'sd32762;
			10'd772:	sine_sample = 16'sd32758;
			10'd773:	sine_sample = 16'sd32753;
			10'd774:	sine_sample = 16'sd32746;
			10'd775:	sine_sample = 16'sd32738;
			10'd776:	sine_sample = 16'sd32729;
			10'd777:	sine_sample = 16'sd32718;
			10'd778:	sine_sample = 16'sd32706;
			10'd779:	sine_sample = 16'sd32693;
			10'd780:	sine_sample = 16'sd32679;
			10'd781:	sine_sample = 16'sd32664;
			10'd782:	sine_sample = 16'sd32647;
			10'd783:	sine_sample = 16'sd32629;
			10'd784:	sine_sample = 16'sd32610;
			10'd785:	sine_sample = 16'sd32590;
			10'd786:	sine_sample = 16'sd32568;
			10'd787:	sine_sample = 16'sd32546;
			10'd788:	sine_sample = 16'sd32522;
			10'd789:	sine_sample = 16'sd32496;
			10'd790:	sine_sample = 16'sd32470;
			10'd791:	sine_sample = 16'sd32442;
			10'd792:	sine_sample = 16'sd32413;
			10'd793:	sine_sample = 16'sd32383;
			10'd794:	sine_sample = 16'sd32352;
			10'd795:	sine_sample = 16'sd32319;
			10'd796:	sine_sample = 16'sd32286;
			10'd797:	sine_sample = 16'sd32251;
			10'd798:	sine_sample = 16'sd32214;
			10'd799:	sine_sample = 16'sd32177;
			10'd800:	sine_sample = 16'sd32138;
			10'd801:	sine_sample = 16'sd32099;
			10'd802:	sine_sample = 16'sd32058;
			10'd803:	sine_sample = 16'sd32015;
			10'd804:	sine_sample = 16'sd31972;
			10'd805:	sine_sample = 16'sd31927;
			10'd806:	sine_sample = 16'sd31881;
			10'd807:	sine_sample = 16'sd31834;
			10'd808:	sine_sample = 16'sd31786;
			10'd809:	sine_sample = 16'sd31737;
			10'd810:	sine_sample = 16'sd31686;
			10'd811:	sine_sample = 16'sd31634;
			10'd812:	sine_sample = 16'sd31581;
			10'd813:	sine_sample = 16'sd31527;
			10'd814:	sine_sample = 16'sd31471;
			10'd815:	sine_sample = 16'sd31415;
			10'd816:	sine_sample = 16'sd31357;
			10'd817:	sine_sample = 16'sd31298;
			10'd818:	sine_sample = 16'sd31238;
			10'd819:	sine_sample = 16'sd31177;
			10'd820:	sine_sample = 16'sd31114;
			10'd821:	sine_sample = 16'sd31050;
			10'd822:	sine_sample = 16'sd30986;
			10'd823:	sine_sample = 16'sd30920;
			10'd824:	sine_sample = 16'sd30853;
			10'd825:	sine_sample = 16'sd30784;
			10'd826:	sine_sample = 16'sd30715;
			10'd827:	sine_sample = 16'sd30644;
			10'd828:	sine_sample = 16'sd30572;
			10'd829:	sine_sample = 16'sd30499;
			10'd830:	sine_sample = 16'sd30425;
			10'd831:	sine_sample = 16'sd30350;
			10'd832:	sine_sample = 16'sd30274;
			10'd833:	sine_sample = 16'sd30196;
			10'd834:	sine_sample = 16'sd30118;
			10'd835:	sine_sample = 16'sd30038;
			10'd836:	sine_sample = 16'sd29957;
			10'd837:	sine_sample = 16'sd29875;
			10'd838:	sine_sample = 16'sd29792;
			10'd839:	sine_sample = 16'sd29707;
			10'd840:	sine_sample = 16'sd29622;
			10'd841:	sine_sample = 16'sd29535;
			10'd842:	sine_sample = 16'sd29448;
			10'd843:	sine_sample = 16'sd29359;
			10'd844:	sine_sample = 16'sd29269;
			10'd845:	sine_sample = 16'sd29178;
			10'd846:	sine_sample = 16'sd29086;
			10'd847:	sine_sample = 16'sd28993;
			10'd848:	sine_sample = 16'sd28899;
			10'd849:	sine_sample = 16'sd28803;
			10'd850:	sine_sample = 16'sd28707;
			10'd851:	sine_sample = 16'sd28610;
			10'd852:	sine_sample = 16'sd28511;
			10'd853:	sine_sample = 16'sd28411;
			10'd854:	sine_sample = 16'sd28311;
			10'd855:	sine_sample = 16'sd28209;
			10'd856:	sine_sample = 16'sd28106;
			10'd857:	sine_sample = 16'sd28002;
			10'd858:	sine_sample = 16'sd27897;
			10'd859:	sine_sample = 16'sd27791;
			10'd860:	sine_sample = 16'sd27684;
			10'd861:	sine_sample = 16'sd27576;
			10'd862:	sine_sample = 16'sd27467;
			10'd863:	sine_sample = 16'sd27357;
			10'd864:	sine_sample = 16'sd27246;
			10'd865:	sine_sample = 16'sd27133;
			10'd866:	sine_sample = 16'sd27020;
			10'd867:	sine_sample = 16'sd26906;
			10'd868:	sine_sample = 16'sd26791;
			10'd869:	sine_sample = 16'sd26674;
			10'd870:	sine_sample = 16'sd26557;
			10'd871:	sine_sample = 16'sd26439;
			10'd872:	sine_sample = 16'sd26320;
			10'd873:	sine_sample = 16'sd26199;
			10'd874:	sine_sample = 16'sd26078;
			10'd875:	sine_sample = 16'sd25956;
			10'd876:	sine_sample = 16'sd25833;
			10'd877:	sine_sample = 16'sd25708;
			10'd878:	sine_sample = 16'sd25583;
			10'd879:	sine_sample = 16'sd25457;
			10'd880:	sine_sample = 16'sd25330;
			10'd881:	sine_sample = 16'sd25202;
			10'd882:	sine_sample = 16'sd25073;
			10'd883:	sine_sample = 16'sd24943;
			10'd884:	sine_sample = 16'sd24812;
			10'd885:	sine_sample = 16'sd24680;
			10'd886:	sine_sample = 16'sd24548;
			10'd887:	sine_sample = 16'sd24414;
			10'd888:	sine_sample = 16'sd24279;
			10'd889:	sine_sample = 16'sd24144;
			10'd890:	sine_sample = 16'sd24008;
			10'd891:	sine_sample = 16'sd23870;
			10'd892:	sine_sample = 16'sd23732;
			10'd893:	sine_sample = 16'sd23593;
			10'd894:	sine_sample = 16'sd23453;
			10'd895:	sine_sample = 16'sd23312;
			10'd896:	sine_sample = 16'sd23170;
			10'd897:	sine_sample = 16'sd23028;
			10'd898:	sine_sample = 16'sd22884;
			10'd899:	sine_sample = 16'sd22740;
			10'd900:	sine_sample = 16'sd22595;
			10'd901:	sine_sample = 16'sd22449;
			10'd902:	sine_sample = 16'sd22302;
			10'd903:	sine_sample = 16'sd22154;
			10'd904:	sine_sample = 16'sd22006;
			10'd905:	sine_sample = 16'sd21856;
			10'd906:	sine_sample = 16'sd21706;
			10'd907:	sine_sample = 16'sd21555;
			10'd908:	sine_sample = 16'sd21403;
			10'd909:	sine_sample = 16'sd21251;
			10'd910:	sine_sample = 16'sd21097;
			10'd911:	sine_sample = 16'sd20943;
			10'd912:	sine_sample = 16'sd20788;
			10'd913:	sine_sample = 16'sd20632;
			10'd914:	sine_sample = 16'sd20475;
			10'd915:	sine_sample = 16'sd20318;
			10'd916:	sine_sample = 16'sd20160;
			10'd917:	sine_sample = 16'sd20001;
			10'd918:	sine_sample = 16'sd19841;
			10'd919:	sine_sample = 16'sd19681;
			10'd920:	sine_sample = 16'sd19520;
			10'd921:	sine_sample = 16'sd19358;
			10'd922:	sine_sample = 16'sd19195;
			10'd923:	sine_sample = 16'sd19032;
			10'd924:	sine_sample = 16'sd18868;
			10'd925:	sine_sample = 16'sd18703;
			10'd926:	sine_sample = 16'sd18538;
			10'd927:	sine_sample = 16'sd18372;
			10'd928:	sine_sample = 16'sd18205;
			10'd929:	sine_sample = 16'sd18037;
			10'd930:	sine_sample = 16'sd17869;
			10'd931:	sine_sample = 16'sd17700;
			10'd932:	sine_sample = 16'sd17531;
			10'd933:	sine_sample = 16'sd17361;
			10'd934:	sine_sample = 16'sd17190;
			10'd935:	sine_sample = 16'sd17018;
			10'd936:	sine_sample = 16'sd16846;
			10'd937:	sine_sample = 16'sd16673;
			10'd938:	sine_sample = 16'sd16500;
			10'd939:	sine_sample = 16'sd16326;
			10'd940:	sine_sample = 16'sd16151;
			10'd941:	sine_sample = 16'sd15976;
			10'd942:	sine_sample = 16'sd15800;
			10'd943:	sine_sample = 16'sd15624;
			10'd944:	sine_sample = 16'sd15447;
			10'd945:	sine_sample = 16'sd15269;
			10'd946:	sine_sample = 16'sd15091;
			10'd947:	sine_sample = 16'sd14912;
			10'd948:	sine_sample = 16'sd14733;
			10'd949:	sine_sample = 16'sd14553;
			10'd950:	sine_sample = 16'sd14373;
			10'd951:	sine_sample = 16'sd14192;
			10'd952:	sine_sample = 16'sd14010;
			10'd953:	sine_sample = 16'sd13828;
			10'd954:	sine_sample = 16'sd13646;
			10'd955:	sine_sample = 16'sd13463;
			10'd956:	sine_sample = 16'sd13279;
			10'd957:	sine_sample = 16'sd13095;
			10'd958:	sine_sample = 16'sd12910;
			10'd959:	sine_sample = 16'sd12725;
			10'd960:	sine_sample = 16'sd12540;
			10'd961:	sine_sample = 16'sd12354;
			10'd962:	sine_sample = 16'sd12167;
			10'd963:	sine_sample = 16'sd11980;
			10'd964:	sine_sample = 16'sd11793;
			10'd965:	sine_sample = 16'sd11605;
			10'd966:	sine_sample = 16'sd11417;
			10'd967:	sine_sample = 16'sd11228;
			10'd968:	sine_sample = 16'sd11039;
			10'd969:	sine_sample = 16'sd10850;
			10'd970:	sine_sample = 16'sd10660;
			10'd971:	sine_sample = 16'sd10469;
			10'd972:	sine_sample = 16'sd10279;
			10'd973:	sine_sample = 16'sd10088;
			10'd974:	sine_sample = 16'sd9896;
			10'd975:	sine_sample = 16'sd9704;
			10'd976:	sine_sample = 16'sd9512;
			10'd977:	sine_sample = 16'sd9319;
			10'd978:	sine_sample = 16'sd9127;
			10'd979:	sine_sample = 16'sd8933;
			10'd980:	sine_sample = 16'sd8740;
			10'd981:	sine_sample = 16'sd8546;
			10'd982:	sine_sample = 16'sd8351;
			10'd983:	sine_sample = 16'sd8157;
			10'd984:	sine_sample = 16'sd7962;
			10'd985:	sine_sample = 16'sd7767;
			10'd986:	sine_sample = 16'sd7571;
			10'd987:	sine_sample = 16'sd7376;
			10'd988:	sine_sample = 16'sd7180;
			10'd989:	sine_sample = 16'sd6983;
			10'd990:	sine_sample = 16'sd6787;
			10'd991:	sine_sample = 16'sd6590;
			10'd992:	sine_sample = 16'sd6393;
			10'd993:	sine_sample = 16'sd6195;
			10'd994:	sine_sample = 16'sd5998;
			10'd995:	sine_sample = 16'sd5800;
			10'd996:	sine_sample = 16'sd5602;
			10'd997:	sine_sample = 16'sd5404;
			10'd998:	sine_sample = 16'sd5205;
			10'd999:	sine_sample = 16'sd5007;
			10'd1000:	sine_sample = 16'sd4808;
			10'd1001:	sine_sample = 16'sd4609;
			10'd1002:	sine_sample = 16'sd4410;
			10'd1003:	sine_sample = 16'sd4211;
			10'd1004:	sine_sample = 16'sd4011;
			10'd1005:	sine_sample = 16'sd3812;
			10'd1006:	sine_sample = 16'sd3612;
			10'd1007:	sine_sample = 16'sd3412;
			10'd1008:	sine_sample = 16'sd3212;
			10'd1009:	sine_sample = 16'sd3012;
			10'd1010:	sine_sample = 16'sd2811;
			10'd1011:	sine_sample = 16'sd2611;
			10'd1012:	sine_sample = 16'sd2411;
			10'd1013:	sine_sample = 16'sd2210;
			10'd1014:	sine_sample = 16'sd2009;
			10'd1015:	sine_sample = 16'sd1809;
			10'd1016:	sine_sample = 16'sd1608;
			10'd1017:	sine_sample = 16'sd1407;
			10'd1018:	sine_sample = 16'sd1206;
			10'd1019:	sine_sample = 16'sd1005;
			10'd1020:	sine_sample = 16'sd804;
			10'd1021:	sine_sample = 16'sd603;
			10'd1022:	sine_sample = 16'sd402;
			10'd1023:	sine_sample = 16'sd201;
			default: sine_sample = 16'sd0;
		endcase
	end
endmodule
