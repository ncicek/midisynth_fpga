module tuning_code_lookup(
	//input wire i_clk,
	input wire [6:0] midi_byte,
	output reg [31:0] tuning_code
);

	always @(midi_byte) begin
		case(midi_byte)
			7'd0:	tuning_code = 32'd1685510;
			7'd1:	tuning_code = 32'd1785736;
			7'd2:	tuning_code = 32'd1891921;
			7'd3:	tuning_code = 32'd2004420;
			7'd4:	tuning_code = 32'd2123609;
			7'd5:	tuning_code = 32'd2249886;
			7'd6:	tuning_code = 32'd2383671;
			7'd7:	tuning_code = 32'd2525411;
			7'd8:	tuning_code = 32'd2675580;
			7'd9:	tuning_code = 32'd2834678;
			7'd10:	tuning_code = 32'd3003237;
			7'd11:	tuning_code = 32'd3181819;
			7'd12:	tuning_code = 32'd3371020;
			7'd13:	tuning_code = 32'd3571471;
			7'd14:	tuning_code = 32'd3783842;
			7'd15:	tuning_code = 32'd4008841;
			7'd16:	tuning_code = 32'd4247219;
			7'd17:	tuning_code = 32'd4499771;
			7'd18:	tuning_code = 32'd4767342;
			7'd19:	tuning_code = 32'd5050823;
			7'd20:	tuning_code = 32'd5351160;
			7'd21:	tuning_code = 32'd5669357;
			7'd22:	tuning_code = 32'd6006474;
			7'd23:	tuning_code = 32'd6363638;
			7'd24:	tuning_code = 32'd6742039;
			7'd25:	tuning_code = 32'd7142942;
			7'd26:	tuning_code = 32'd7567683;
			7'd27:	tuning_code = 32'd8017681;
			7'd28:	tuning_code = 32'd8494437;
			7'd29:	tuning_code = 32'd8999543;
			7'd30:	tuning_code = 32'd9534684;
			7'd31:	tuning_code = 32'd10101645;
			7'd32:	tuning_code = 32'd10702321;
			7'd33:	tuning_code = 32'd11338714;
			7'd34:	tuning_code = 32'd12012949;
			7'd35:	tuning_code = 32'd12727276;
			7'd36:	tuning_code = 32'd13484079;
			7'd37:	tuning_code = 32'd14285884;
			7'd38:	tuning_code = 32'd15135367;
			7'd39:	tuning_code = 32'd16035363;
			7'd40:	tuning_code = 32'd16988875;
			7'd41:	tuning_code = 32'd17999086;
			7'd42:	tuning_code = 32'd19069367;
			7'd43:	tuning_code = 32'd20203291;
			7'd44:	tuning_code = 32'd21404641;
			7'd45:	tuning_code = 32'd22677427;
			7'd46:	tuning_code = 32'd24025897;
			7'd47:	tuning_code = 32'd25454552;
			7'd48:	tuning_code = 32'd26968158;
			7'd49:	tuning_code = 32'd28571768;
			7'd50:	tuning_code = 32'd30270734;
			7'd51:	tuning_code = 32'd32070725;
			7'd52:	tuning_code = 32'd33977750;
			7'd53:	tuning_code = 32'd35998172;
			7'd54:	tuning_code = 32'd38138735;
			7'd55:	tuning_code = 32'd40406582;
			7'd56:	tuning_code = 32'd42809282;
			7'd57:	tuning_code = 32'd45354855;
			7'd58:	tuning_code = 32'd48051795;
			7'd59:	tuning_code = 32'd50909103;
			7'd60:	tuning_code = 32'd53936316;
			7'd61:	tuning_code = 32'd57143536;
			7'd62:	tuning_code = 32'd60541468;
			7'd63:	tuning_code = 32'd64141451;
			7'd64:	tuning_code = 32'd67955500;
			7'd65:	tuning_code = 32'd71996344;
			7'd66:	tuning_code = 32'd76277469;
			7'd67:	tuning_code = 32'd80813164;
			7'd68:	tuning_code = 32'd85618565;
			7'd69:	tuning_code = 32'd90709709;
			7'd70:	tuning_code = 32'd96103589;
			7'd71:	tuning_code = 32'd101818206;
			7'd72:	tuning_code = 32'd107872632;
			7'd73:	tuning_code = 32'd114287072;
			7'd74:	tuning_code = 32'd121082935;
			7'd75:	tuning_code = 32'd128282901;
			7'd76:	tuning_code = 32'd135910999;
			7'd77:	tuning_code = 32'd143992688;
			7'd78:	tuning_code = 32'd152554939;
			7'd79:	tuning_code = 32'd161626327;
			7'd80:	tuning_code = 32'd171237129;
			7'd81:	tuning_code = 32'd181419419;
			7'd82:	tuning_code = 32'd192207179;
			7'd83:	tuning_code = 32'd203636412;
			7'd84:	tuning_code = 32'd215745263;
			7'd85:	tuning_code = 32'd228574144;
			7'd86:	tuning_code = 32'd242165870;
			7'd87:	tuning_code = 32'd256565802;
			7'd88:	tuning_code = 32'd271821999;
			7'd89:	tuning_code = 32'd287985376;
			7'd90:	tuning_code = 32'd305109877;
			7'd91:	tuning_code = 32'd323252655;
			7'd92:	tuning_code = 32'd342474258;
			7'd93:	tuning_code = 32'd362838837;
			7'd94:	tuning_code = 32'd384414357;
			7'd95:	tuning_code = 32'd407272824;
			7'd96:	tuning_code = 32'd431490527;
			7'd97:	tuning_code = 32'd457148289;
			7'd98:	tuning_code = 32'd484331740;
			7'd99:	tuning_code = 32'd513131604;
			7'd100:	tuning_code = 32'd543643997;
			7'd101:	tuning_code = 32'd575970752;
			7'd102:	tuning_code = 32'd610219755;
			7'd103:	tuning_code = 32'd646505310;
			7'd104:	tuning_code = 32'd684948516;
			7'd105:	tuning_code = 32'd725677674;
			7'd106:	tuning_code = 32'd768828714;
			7'd107:	tuning_code = 32'd814545649;
			7'd108:	tuning_code = 32'd862981054;
			7'd109:	tuning_code = 32'd914296577;
			7'd110:	tuning_code = 32'd968663481;
			7'd111:	tuning_code = 32'd1026263209;
			7'd112:	tuning_code = 32'd1087287995;
			7'd113:	tuning_code = 32'd1151941504;
			7'd114:	tuning_code = 32'd1220439510;
			7'd115:	tuning_code = 32'd1293010620;
			7'd116:	tuning_code = 32'd1369897032;
			7'd117:	tuning_code = 32'd1451355349;
			7'd118:	tuning_code = 32'd1537657429;
			7'd119:	tuning_code = 32'd1629091297;
			7'd120:	tuning_code = 32'd1725962107;
			7'd121:	tuning_code = 32'd1828593155;
			7'd122:	tuning_code = 32'd1937326962;
			7'd123:	tuning_code = 32'd2052526418;
			7'd124:	tuning_code = 32'd2174575990;
			7'd125:	tuning_code = 32'd2303883007;
			7'd126:	tuning_code = 32'd2440879020;
			7'd127:	tuning_code = 32'd2586021239;

			default: tuning_code <= 32'd66213;
		endcase
	end
endmodule
